`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Project: Bubble Sort
// Module Name:Incrementer
//////////////////////////////////////////////////////////////////////////////////
module dp_inc(a,b);
parameter  datawidth = 8;
input [datawidth-1:0] a;
output reg [datawidth-1:0] b;

always@(a) begin
	b<=a+1;
end


endmodule
